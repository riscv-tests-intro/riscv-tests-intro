package miriscv_test_pkg;

  `include "mem_model.sv"
  `include "miriscv_mem_item.sv"
  `include "miriscv_mem_seq.sv"
  `include "miriscv_mem_monitor.sv"
  `include "miriscv_mem_driver.sv"
  `include "miriscv_mem_agent.sv"
  `include "miriscv_rvfi_item.sv"
  `include "miriscv_rvfi_monitor.sv"
  `include "miriscv_hammer_dpi.svh"
  `include "miriscv_scoreboard.sv"
  `include "miriscv_test.sv"

endpackage