typedef struct {
    bit [31:0] pc;
    bit [31:0] bits;
    bit [31:0] rd;
    string     str;
} miriscv_insn_info_s;
